------------------------------------------------------------------------------------------------
--
--  DISTRIBUTED HEMPS  - version 5.0
--
--  Research group: GAPH-PUCRS    -    contact   fernando.moraes@pucrs.br
--
--  Distribution:  November 2015
--
--  Source name:  seek_pkg.vhd
--
--  Brief description:  Functions and constants for seek module.
--
------------------------------------------------------------------------------------------------

library IEEE;
use IEEE.Std_Logic_1164.all;
use IEEE.std_logic_unsigned.all;
use work.standards.all;

package seek_pkg is

	constant	NPORT_SEEK								: integer := 5;
	--WARNING : modify source target size to 8
	constant	TARGET_SIZE								: integer := 16;
	constant	SOURCE_SIZE								: integer := 32;
	constant	SEEK_PAYLOAD_SIZE						: integer := 8;
	constant	TAM_SERVICE_SEEK						: integer := 6;

	constant	EAST									: integer := 0;
	constant	WEST									: integer := 1;
	constant	NORTH									: integer := 2;
	constant	SOUTH									: integer := 3;
	constant	LOCAL									: integer := 4;

	constant	ROW0									: integer := 0;
	constant	ROW1									: integer := 1;
	constant	ROW2									: integer := 2;
	constant	ROW3									: integer := 3;
	constant	ROW4									: integer := 4;
	constant	ROW5									: integer := 5;
	constant	ROW6									: integer := 6;
	constant	ROW7									: integer := 7;

--table sizes
    constant    TABLE_HEIGHT							: integer := 8;
    constant    TABLE_SEEK_LENGHT						: integer := 8;
-- ordem SET_SECURE_ZONE_SERVICE, SET_EXCESS_SZ_SERVICE, SECURE_ZONE_CLOSED_SERVICE
-- OPEN_SECURE_ZONE_SERVICE, SECURE_ZONE_OPENED_SERVICE
-- PDN services
    constant    START_APP_SERVICE                       : std_logic_vector(TAM_SERVICE_SEEK-1 downto 0) := "000001";
    constant    TARGET_UNREACHABLE_SERVICE              : std_logic_vector(TAM_SERVICE_SEEK-1 downto 0) := "000010";
    constant    CLEAR_SERVICE                           : std_logic_vector(TAM_SERVICE_SEEK-1 downto 0) := "000011";
    constant    BACKTRACK_SERVICE                       : std_logic_vector(TAM_SERVICE_SEEK-1 downto 0) := "000100";
    constant    SEARCHPATH_SERVICE                      : std_logic_vector(TAM_SERVICE_SEEK-1 downto 0) := "000101";
    constant    END_TASK_SERVICE                        : std_logic_vector(TAM_SERVICE_SEEK-1 downto 0) := "000110";
    constant    SET_SECURE_ZONE_SERVICE                 : std_logic_vector(TAM_SERVICE_SEEK-1 downto 0) := "000111";
    constant    PACKET_RESEND_SERVICE                   : std_logic_vector(TAM_SERVICE_SEEK-1 downto 0) := "001000";
    constant    WARD_SERVICE                            : std_logic_vector(TAM_SERVICE_SEEK-1 downto 0) := "001001";
    constant    OPEN_SECURE_ZONE_SERVICE                : std_logic_vector(TAM_SERVICE_SEEK-1 downto 0) := "001010";
    constant    SECURE_ZONE_CLOSED_SERVICE              : std_logic_vector(TAM_SERVICE_SEEK-1 downto 0) := "001011";
    constant    SECURE_ZONE_OPENED_SERVICE              : std_logic_vector(TAM_SERVICE_SEEK-1 downto 0) := "001100";
    constant    FREEZE_TASK_SERVICE                     : std_logic_vector(TAM_SERVICE_SEEK-1 downto 0) := "001101";
    constant    UNFREEZE_TASK_SERVICE                   : std_logic_vector(TAM_SERVICE_SEEK-1 downto 0) := "001110";
    constant    MASTER_CANDIDATE_SERVICE                : std_logic_vector(TAM_SERVICE_SEEK-1 downto 0) := "001111";
    constant    TASK_ALLOCATED_SERVICE                  : std_logic_vector(TAM_SERVICE_SEEK-1 downto 0) := "010000";
    constant    INITIALIZE_SLAVE_SERVICE                : std_logic_vector(TAM_SERVICE_SEEK-1 downto 0) := "010001";
    constant    INITIALIZE_CLUSTER_SERVICE              : std_logic_vector(TAM_SERVICE_SEEK-1 downto 0) := "010010";
    constant    LOAN_PROCESSOR_REQUEST_SERVICE          : std_logic_vector(TAM_SERVICE_SEEK-1 downto 0) := "010011"; --
    constant    LOAN_PROCESSOR_RELEASE_SERVICE          : std_logic_vector(TAM_SERVICE_SEEK-1 downto 0) := "010100"; --
    constant    END_TASK_OTHER_CLUSTER_SERVICE          : std_logic_vector(TAM_SERVICE_SEEK-1 downto 0) := "010101";
    constant    WAIT_KERNEL_SERVICE                     : std_logic_vector(TAM_SERVICE_SEEK-1 downto 0) := "010110";
    constant    SEND_KERNEL_SERVICE                     : std_logic_vector(TAM_SERVICE_SEEK-1 downto 0) := "010111";
    constant    WAIT_KERNEL_SERVICE_ACK                 : std_logic_vector(TAM_SERVICE_SEEK-1 downto 0) := "011000";
    constant    FAIL_KERNEL_SERVICE                     : std_logic_vector(TAM_SERVICE_SEEK-1 downto 0) := "011001";
    constant    NEW_APP_SERVICE                         : std_logic_vector(TAM_SERVICE_SEEK-1 downto 0) := "011010";
    constant    NEW_APP_ACK_SERVICE                     : std_logic_vector(TAM_SERVICE_SEEK-1 downto 0) := "011011";
    constant    GMV_READY_SERVICE                       : std_logic_vector(TAM_SERVICE_SEEK-1 downto 0) := "011100";
    constant    SET_SZ_RECEIVED_SERVICE                 : std_logic_vector(TAM_SERVICE_SEEK-1 downto 0) := "011101";
    constant    SET_EXCESS_SZ_SERVICE                   : std_logic_vector(TAM_SERVICE_SEEK-1 downto 0) := "011110";
    constant    RCV_FREEZE_TASK_SERVICE                 : std_logic_vector(TAM_SERVICE_SEEK-1 downto 0) := "011111";
    constant    BR_TO_APPID_SERVICE                     : std_logic_vector(TAM_SERVICE_SEEK-1 downto 0) := "100000";
    constant    SET_AP_SERVICE                          : std_logic_vector(TAM_SERVICE_SEEK-1 downto 0) := "100001";
    constant    MSG_DELIVERY_CONTROL                    : std_logic_vector(TAM_SERVICE_SEEK-1 downto 0) := "100010";
    constant    MSG_REQUEST_CONTROL                     : std_logic_vector(TAM_SERVICE_SEEK-1 downto 0) := "100011";
    constant    RENEW_KEY                               : std_logic_vector(TAM_SERVICE_SEEK-1 downto 0) := "100100";
    constant    KEY_ACK                                 : std_logic_vector(TAM_SERVICE_SEEK-1 downto 0) := "100101";
    constant    REQUEST_SNIP_RENEWAL                    : std_logic_vector(TAM_SERVICE_SEEK-1 downto 0) := "100110";
    constant    LC_NOTIFICATION                         : std_logic_vector(TAM_SERVICE_SEEK-1 downto 0) := "100111";
    constant    AP_NOTIFICATION                         : std_logic_vector(TAM_SERVICE_SEEK-1 downto 0) := "101000";
    constant    UNEXPECTED_DATA                         : std_logic_vector(TAM_SERVICE_SEEK-1 downto 0) := "101001";
    constant    MISSING_PACKET                          : std_logic_vector(TAM_SERVICE_SEEK-1 downto 0) := "101010";
    constant    PROBE_REQUEST                           : std_logic_vector(TAM_SERVICE_SEEK-1 downto 0) := "101011";
    constant    PROBE_PATH                              : std_logic_vector(TAM_SERVICE_SEEK-1 downto 0) := "101100";
    constant    PROBE_CONTROL                           : std_logic_vector(TAM_SERVICE_SEEK-1 downto 0) := "101101";
    constant    PROBE_RESULT                            : std_logic_vector(TAM_SERVICE_SEEK-1 downto 0) := "101110";
    constant    PROBE_REQUEST_PATH                      : std_logic_vector(TAM_SERVICE_SEEK-1 downto 0) := "101111";
    constant    PROBE_PATH_XY                           : std_logic_vector(TAM_SERVICE_SEEK-1 downto 0) := "110000";
    constant    RESET_HERMES_PORT_SERVICE               : std_logic_vector(TAM_SERVICE_SEEK-1 downto 0) := "110001";
    constant    INIT_ROUTER_RESET                       : std_logic_vector(TAM_SERVICE_SEEK-1 downto 0) := "110010";
    constant    REPORT_SUSPICIOUS_PATH                  : std_logic_vector(TAM_SERVICE_SEEK-1 downto 0) := "110011";

	subtype		regNtarget								is std_logic_vector((TARGET_SIZE-1) downto 0);
	subtype		regNsource								is std_logic_vector((SOURCE_SIZE-1) downto 0);
	subtype		regNpayload								is std_logic_vector((SEEK_PAYLOAD_SIZE-1) downto 0);

	type		regNportNsource_neighbor				is array (0 to NPORT_SEEK-1) of regNsource;
	type		regNportNtarget_neighbor				is array (0 to NPORT_SEEK-1) of regNtarget;
	type		regNportNpayload_neighbor				is array (0 to NPORT_SEEK-1) of regNpayload;

    subtype     seek_bitN_service                       is std_logic_vector(TAM_SERVICE_SEEK-1 downto 0);
    type        regNport_seek_bitN_service              is array (NPORT_SEEK-1 downto 0) of seek_bitN_service;
	
    constant	REG_BACKTRACK_SIZE						: integer := 96;

    -- table
	type		source_table_type						is array (TABLE_SEEK_LENGHT-1 downto 0) of regNsource;
	type		target_table_type						is array (TABLE_SEEK_LENGHT-1 downto 0) of regNtarget;
	type		service_table_type						is array (TABLE_SEEK_LENGHT-1 downto 0) of seek_bitN_service;
	type		payload_table_type						is array (TABLE_SEEK_LENGHT-1 downto 0) of regNpayload;
	type		backtrack_port_table_type 				is array (TABLE_SEEK_LENGHT-1 downto 0) of std_logic_vector(2 downto 0);
	type		source_router_port_table_type			is array (TABLE_SEEK_LENGHT-1 downto 0) of std_logic_vector(1 downto 0);

	-- output FSM States

	type T_ea_manager is (S_INIT, ARBITRATION, TEST_SERVICE, SERVICE_BACKTRACK, BACKTRACK_PROPAGATE, INIT_BACKTRACK, PREPARE_NEXT,
		BACKTRACK_MOUNT, CLEAR_TABLE, COMPARE_TARGET, SEND_LOCAL, PROPAGATE, WAIT_ACK_PORTS, INIT_CLEAR, END_BACKTRACK, COUNT, HERMES_RESET);
	
	-- input FSM States

	type T_ea_manager_input is (S_INIT_INPUT, ARBITRATION_INPUT, LOOK_TABLE_INPUT, TEST_SPACE_AVAIL, SERVICE_INPUT, TABLE_WRITE_INPUT,
		WRITE_BACKTRACK_INPUT, TEST_SEND_LOCAL, WRITE_CLEAR_INPUT, WAIT_REQ_DOWN, WAIT_REQ_DOWN_NACK, SEND_NACK);


end package seek_pkg;

----------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- Service                      type                        	Operation Mode      Payload     Target                          Source
-- START_APP_SERVICE            Broadcast to all local ports   	Global              AppID       RH_corner                       --
-- TARGET_UNREACHABLE_SERVICE   Broadcast With Target       	Global              --          TaskID Address                  --
-- CLEAR_SERVICE                Broadcast Without Target    	Global              --          --                              --
-- BACKTRACK_SERVICE            Unicast                     	Restrict            Hop number  --                              --
-- SEARCHPATH_SERVICE           Broadcast With Target          	Restrict            Hop number  Target Unreachable Address
-- END_TASK_SERVICE             Broadcast With Target       	Global              TaskID      CMP Address
-- PACKET_RESEND_SERVICE        Broadcast With Target       	Global              --          TaskID Address
-- WARD_SERVICE                 Broadcast With Target       	Global              --          CMP WARD Address
-- SET_SECURE_ZONE              Broadcast to all local ports    Global              RH_corner   LL_corner
-- OPEN_SECURE_ZONE             Broadcast to all local ports    Global              RH_corner   AppID
-- SECURE_ZONE_CLOSED           Broadcast With Target           Global              RH_corner   CMP Address -- cluster manager pe (target)
-- SECURE_ZONE_OPENED           Broadcast With Target           Global              AppID       CMP Address
-- FREEZE_TASK_SERVICE          Broadcast to all local ports    Global              0           CMP WARD Address
-- UNFREEZE_TASK_SERVICE        Broadcast to all local ports    Global              0           CMP WARD Address
-- MASTER_CANDIDATE_SERVICE     Broadcast With Target           Global              0           CMP WARD Address
-- TASK_ALLOCATED_SERVICE       Broadcast With Target           Global              TaskID      CMP Address
-- INITIALIZE_SLAVE_SERVICE     Broadcast to all local ports    Global              RH_corner   LL_corner
-- WAIT_KERNEL_SERVICE          Broadcast With Target           Global              ?           Next master of cluster
-- SEND_KERNEL_SERVICE          Broadcast With Target           Global              ?           Master fail of cluster
-- FAIL_KERNEL_SERVICE          Broadcast With Target           Global              ?           CMP WARD Address
-- NEW_APP_SERVICE              Broadcast to all local ports    Global              Nr,task     Global master virtual
-- NEW_APP_ACK_SERVICE          Broadcast With Target           Global              Nr,task     Address of the LMP
-- GMV_READY_SERVICE            Broadcast Without Target        Global              --          Injection Entity 
-- MSG_DELIVERY_CONTROL             Broadcast With Target           Global              TgtAppID    TargetID                        SrcAppID
-- MSG_REQUEST_CONTROL          Broadcast With Target           Global              TgtAppID    TargetID                        SrcAppID

--Seek(MSG_DELIVERY_CONTROL, target, (AppID << 16), 0); 
